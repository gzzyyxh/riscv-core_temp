`include "defines.v"

module ctrl(

	input wire										rst,
	
	input wire							stallreq_from_if,
	input wire							stallreq_from_mem,

	input wire                   stallreq_from_id,

  //来自执行阶段的暂停请求
	input wire                   stallreq_from_ex,
	
	input wire[31:0]					excepttype_i,
	input wire[`RegBus]				csr_mepc_i,
	input wire[`RegBus]				csr_mtvec_i,
	
	output reg[5:0]              stall,
	
	output reg[`RegBus]				new_pc,
	output reg							flush
	
);


	always @ (*) begin
		if(rst == `RstEnable) begin
			stall <= 6'b000000;
			flush <= 1'b0;
			new_pc <= `ZeroWord;
		end else if(excepttype_i != `ZeroWord) begin
			flush <= 1'b1;
			stall <= 6'b000000;
			case(excepttype_i)
				32'h00000001:		begin
//					new_pc <= {csr_mtvec_i[31:2], 2'b00};		//??????????????
					new_pc <= 32'h00000020;
				end
				32'h00000008, 32'h0000000a:		begin
//					new_pc <= {csr_mtvec_i[31:2], 2'b00};		//??????????????
					new_pc <= 32'h00000040;
				end
				32'h0000000e:		begin
					new_pc <= csr_mepc_i;
				end
				default:		begin
				end
			endcase
		end else if(stallreq_from_mem == `Stop) begin
			stall <= 6'b011111;
			flush <= 1'b0;
		end else if(stallreq_from_ex == `Stop) begin
			stall <= 6'b001111;
			flush <= 1'b0;
		end else if(stallreq_from_id == `Stop) begin
			stall <= 6'b000111;		
			flush <= 1'b0;
		end else if(stallreq_from_if == `Stop) begin
			stall <= 6'b000011;										//忽略延迟槽
			flush <= 1'b0;
		end else begin
			stall <= 6'b000000;
			flush <= 1'b0;
			new_pc <= `ZeroWord;
		end    //if
	end      //always
			

endmodule